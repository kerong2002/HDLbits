//2022_11_9 kerong
//Serial receiver and datapath
module top_module(
    input clk,
    input in,
    input reset,    // Synchronous reset
    output [7:0] out_byte,
    output done
); //
    

    // Use FSM from Fsm_serial

    // New: Datapath to latch input bits.

endmodule
