//2022_11_9 kerong
//One-hot FSM
module top_module(
    input in,
    input [9:0] state,
    output [9:0] next_state,
    output out1,
    output out2);

endmodule
