//2022/09/22 陳科融
//GND
module top_module (
    output out);

assign out = 1'b0;

endmodule
