//2022-02-22 陳科融
//Simple wire
module top_module( input in, output out );

assign  out=in;

endmodule