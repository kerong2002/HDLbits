//2022_11_10 kerong
//Combinational circuit 1
module top_module (
    input a,
    input b,
    output q );//

    assign q = a & b; // Fix me

endmodule
