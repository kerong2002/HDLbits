//2022-02-22 陳科融
//Getting start
module top_module( output one );

// Insert your code here
    assign one = 1'b1;

endmodule
