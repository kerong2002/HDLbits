//2022-09/22 陳科融
//Wire
module top_module (
    input in,
    output out);

assign  out = in;

endmodule
