//2022-02-22 陳科融
//Output zero
module top_module(
    output zero
);// Module body starts after semicolon

assign zero=0;

endmodule
