//2022_11_1 kerong
//3-variable
module top_module(
    input a,
    input b,
    input c,
    output out  ); 

assign out = a | b | c;

endmodule
